'timescale 1ms/100ns
module fsm_vending_machine_tb();
  reg clk,rst,
  reg [1:0]coin,
  wire x,

  
